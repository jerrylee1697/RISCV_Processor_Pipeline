`timescale 1ns / 1ps

module tb_top;

//clock and reset signal declaration
  logic tb_clk, reset;
  logic [31:0] tb_ALU_Result;

    //clock generation
  always #10 tb_clk = ~tb_clk;

  //reset Generation
  initial begin
    tb_clk = 0;
    reset = 1;
    #25 reset =0;
  end


  riscv riscV(
      .clk(tb_clk),
      .reset(reset),
      .WB_Data(tb_ALU_Result)      
     );

  initial begin
    #2000;
    $finish;
   end
endmodule
