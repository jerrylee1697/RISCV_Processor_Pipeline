`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 01/07/2018 10:10:33 PM
// Design Name:
// Module Name: Controller
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module Controller(

    //Input
    input logic [6:0] Opcode, //7-bit opcode field from the instruction

    //Outputs
    output logic ALUSrc,//0: The second ALU operand comes from the second register file output (Read data 2);
                  //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic [1:0]  MemtoReg, //0: The value fed to the register Write data input comes from the ALU.
                     //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic Branch,  //0: branch is not taken; 1: branch is taken
    output logic jalr,
    output logic lui,
    output logic jal,
    output logic ReadFlag,
    output logic WriteFlag,
    output logic [1:0] ALUOp
);

//    localparam R_TYPE = 7'b0110011;
//    localparam LW     = 7'b0000011;
//    localparam SW     = 7'b0100011;
////    localparam BR     = 7'b1100011;
//    localparam RTypeI = 7'b0010011; //addi,ori,andi

    logic [6:0] R_TYPE, LW, SW, RTypeI, JALR, BR, LUI, AUIPC, JAL;

    assign R_TYPE = 7'b0110011;
    assign RTypeI = 7'b0010011; //addi,ori,andi
    assign LW     = 7'b0000011;
    assign SW     = 7'b0100011;
    assign JALR   = 7'b1100111;
    assign BR     = 7'b1100011;
    assign LUI    = 7'b0110111;
    assign AUIPC  = 7'b0010111;
    assign JAL    = 7'b1101111;

  assign ALUSrc   = (Opcode==LW || Opcode==SW || Opcode==RTypeI || Opcode==LUI || Opcode==AUIPC);

  assign MemtoReg = (Opcode==R_TYPE || Opcode==RTypeI) ? 2'b00 :
                    (Opcode==LW) ? 2'b01 :
                    (Opcode==JAL || Opcode==JALR) ? 2'b10 :
                    (Opcode==AUIPC) ? 2'b11 :
                    2'b00;

  assign RegWrite = (Opcode==R_TYPE || Opcode==LW || Opcode == RTypeI || Opcode==JALR || Opcode==JAL || Opcode==AUIPC);
  assign MemRead  = (Opcode==LW);
  assign MemWrite = (Opcode==SW || Opcode==JAL || Opcode==JALR || Opcode==AUIPC);
  assign Branch = (Opcode==BR);
  assign jalr = (Opcode==JALR);
  assign ReadFlag = (Opcode==LW);
  assign WriteFlag = (Opcode==SW);
  //assign ALUOp[0] = 0;
  //assign ALUOp[1] = (Opcode==R_TYPE);
  assign ALUOp[1:0] = (Opcode == R_TYPE) ? 2'b10 :
                      (Opcode == RTypeI) ? 2'b10 :
                      (Opcode == LW)     ? 2'b00 :
                      (Opcode == SW)     ? 2'b00 :
                      (Opcode == JALR)   ? 2'b00 :
                      (Opcode == BR)     ? 2'b01 :
                      (Opcode == LUI)    ? 2'b11 :
                      (Opcode == AUIPC)  ? 2'b11 :
                      (Opcode == JAL)    ? 2'b11 :
                      2'b00;
  assign jal = (Opcode == JAL);
  assign auipc = (Opcode == AUIPC);
  assign lui = (Opcode == LUI);



endmodule

//           Opcode     ALUop
// R-type    0110011    10      Adder
// R-typeI   0010011    10

// Lw        0000011    00      Arithmetic
// Sw        0100011    00
// JALR      1100111    00

// SB        1100011    01  (branches) Adder

// LUI       0110111    11      Comparator
// AUIPC     0010111    11
// JAL       1101111    11
